module datapath (
    clk, reset, RegWrite, ALUSrc, PCSrc, ResultSrc, Jump, fp_RegWrite, add_sub,
    fp_ALUCtrl, Instr, ALUCtrl, ImmSrc, ReadData, PC, ALUResult, WriteData, Zero
);
    input clk, reset, RegWrite, ALUSrc, PCSrc, Jump, fp_RegWrite, add_sub;
    input [1:0] ResultSrc;
    input [31:0] Instr;
    input [1:0] ALUCtrl, ImmSrc;
    input [31:0] ReadData;
    input [3:0] fp_ALUCtrl;
    output wire [31:0] PC;
    output wire [31:0] ALUResult;
    output wire [31:0] WriteData;
    output wire Zero;
    //////////////////////////////////////////////////////////////////////////////////////////
    wire [31:0] RD1, RD2, WD3, PCTarget, PCPlus4, PCNext, ImmExt, TmpResult;
    wire [31:0] TmpResultORfp_ALUResult, TmpPC;
    wire [31:0] fp_RD1, fp_RD2, neg_fp_RD2, fp_WD3, fp_Op1, fp_Op2, fp_ALUResult, fp_ALUResultORReadData;
    wire fp_sw;
    wire [31:0] SrcB;
    //////////////////////////////////////////////////////////////////////////////////////////
    assign neg_fp_RD2 = {~fp_RD2[31] , fp_RD2[30:0]};
    assign fp_sw = Instr[2];
    //Instantiate building blocks 
    add_by_4 add_by_4 (.PC(PC), .PCPlus4(PCPlus4));
    //////////////////////////////////////////////////////////////////////////////////////////
    add_to_ImmExt add_to_ImmExt (PC, ImmExt, TmpPC);
    //////////////////////////////////////////////////////////////////////////////////////////
    PC pc (.clk(clk), .reset(reset), .PC(PC), .PCNext(PCNext));
    //////////////////////////////////////////////////////////////////////////////////////////
    reg_file reg_file (.A1(Instr[19:15]), .A2(Instr[24:20]), .A3(Instr[11:7]),
                        .WE3(RegWrite), .RD1(RD1), .RD2(RD2), .WD3(WD3), .clk(clk));
    //////////////////////////////////////////////////////////////////////////////////////////
    mux_2 i7 (fp_RD1, RD1, & fp_ALUCtrl, fp_Op1);
    //////////////////////////////////////////////////////////////////////////////////////////
    mux_2 i9 (fp_RD2, neg_fp_RD2, add_sub, fp_Op2);
    //////////////////////////////////////////////////////////////////////////////////////////
    fp_alu fp_alu (.A(fp_Op1), .B(fp_Op2), .ALUCtrl(fp_ALUCtrl), .ALUResult(fp_ALUResult));
    //////////////////////////////////////////////////////////////////////////////////////////
    mux_2 i0 (fp_ALUResult, ReadData, ALUSrc, fp_WD3);
    //////////////////////////////////////////////////////////////////////////////////////////
    reg_file fp_reg_file (.A1(Instr[19:15]), .A2(Instr[24:20]), .A3(Instr[11:7]),
                        .WE3(fp_RegWrite), .RD1(fp_RD1), .RD2(fp_RD2), .WD3(fp_WD3), .clk(clk));
    //////////////////////////////////////////////////////////////////////////////////////////
    mux_2 i8 (RD2, fp_RD2, fp_sw, WriteData);
    //////////////////////////////////////////////////////////////////////////////////////////
    imm_ext imm_ext (Instr[31:7], ImmSrc, ImmExt);
    //////////////////////////////////////////////////////////////////////////////////////////
    mux_2 i1 (RD2, ImmExt, ALUSrc, SrcB);
    //////////////////////////////////////////////////////////////////////////////////////////
    alu alu (.A(RD1), .B(SrcB), .ALUCtrl(ALUCtrl), .ALUResult(ALUResult), .Zero(Zero));
    //////////////////////////////////////////////////////////////////////////////////////////
    mux_2 i2 (ALUResult, ReadData, ResultSrc[0], TmpResult);
    //////////////////////////////////////////////////////////////////////////////////////////
    mux_2 i3 (TmpResult, fp_ALUResult, ResultSrc[1], TmpResultORfp_ALUResult);
    //////////////////////////////////////////////////////////////////////////////////////////
    mux_2 i4 (TmpResultORfp_ALUResult, PCPlus4, Jump, WD3);
    //////////////////////////////////////////////////////////////////////////////////////////
    mux_2 i5 (TmpPC, ALUResult, (Jump & ALUSrc), PCTarget);
    //////////////////////////////////////////////////////////////////////////////////////////
    mux_2 i6 (PCPlus4, PCTarget, PCSrc, PCNext);
    //////////////////////////////////////////////////////////////////////////////////////////
    
endmodule