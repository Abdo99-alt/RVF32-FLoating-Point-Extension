localparam N_INF        = 0;
localparam N_NORMAL     = 1;
localparam N_SUBNORMAL  = 2;
localparam N_ZERO       = 3;
localparam ZERO         = 4;
localparam SUBNORMAL    = 5;
localparam NORMAL       = 6;
localparam INF          = 7;
localparam SNAN         = 8;
localparam QNAN         = 9;

localparam NTYPES       = 10;
localparam NEXCEPTIONS  = 5;

localparam EMAX         = 127;
localparam EMIN         = -126;
localparam BIAS         = 127;
localparam NEXP         = 8;
localparam NSIG         = 23;