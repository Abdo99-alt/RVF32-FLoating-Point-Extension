module top (
    clk, reset
);
    input clk, reset;
    //////////////////////////////////////////////////////////////////////////////////////////////////
    wire [31:0] Instr, PC;
    wire [31:0] ALUResult, ReadData, WriteData;
    wire RegWrite, Zero, MemWrite, ALUSrc, PCSrc, Jump, fp_RegWrite, add_sub;
    wire [1:0] ImmSrc, ALUCtrl, ResultSrc;
    wire [3:0] fp_ALUCtrl;
    //////////////////////////////////////////////////////////////////////////////////////////////////
    datapath datapath (clk, reset, RegWrite, ALUSrc, PCSrc, ResultSrc, Jump, fp_RegWrite, add_sub, 
                        fp_ALUCtrl, Instr, ALUCtrl, ImmSrc, ReadData, PC, ALUResult, WriteData, Zero);
    //////////////////////////////////////////////////////////////////////////////////////////////////
    ctrl_unit ctrl_unit (Instr[6:0], Instr[31:27], Instr[14:12], Instr[30], Zero, ImmSrc, ALUCtrl, 
                        RegWrite, ALUSrc, MemWrite, ResultSrc, PCSrc, Jump, fp_RegWrite, add_sub, fp_ALUCtrl);
    //////////////////////////////////////////////////////////////////////////////////////////////////
    instr_mem instr_mem (PC, Instr);
    //////////////////////////////////////////////////////////////////////////////////////////////////
    data_mem data_mem (clk, MemWrite, WriteData, ALUResult, ReadData);
    //////////////////////////////////////////////////////////////////////////////////////////////////
endmodule