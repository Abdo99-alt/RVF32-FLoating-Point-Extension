module fp_cvt(i, f);
    input wire signed [31:0] i;
    output wire [31:0] f;
    ///////////////////////////////////////////////////////////////////
    reg [7:0] fExp;
    reg [4:0] sa;
    reg [30:0] tSig; 
    reg [24:0] roSig;
    reg [31:0] i_unsigned;
    ///////////////////////////////////////////////////////////////////
    always @(*) begin
        if (i[31] == 1'b1) begin
            i_unsigned = (~i) + 1;
        end
        else begin
            i_unsigned = i;
        end
    end
    ///////////////////////////////////////////////////////////////////
    always @(i_unsigned) begin
        casez (i_unsigned)
            32'b01??????????????????????????????: sa = 5'd30;
            32'b001?????????????????????????????: sa = 5'd29;
            32'b0001????????????????????????????: sa = 5'd28;
            32'b00001???????????????????????????: sa = 5'd27;
            32'b000001??????????????????????????: sa = 5'd26;
            32'b0000001?????????????????????????: sa = 5'd25;
            32'b00000001????????????????????????: sa = 5'd24;
            32'b000000001???????????????????????: sa = 5'd23;
            32'b0000000001??????????????????????: sa = 5'd22;
            32'b00000000001?????????????????????: sa = 5'd21;
            32'b000000000001????????????????????: sa = 5'd20;
            32'b0000000000001???????????????????: sa = 5'd19;
            32'b00000000000001??????????????????: sa = 5'd18;
            32'b000000000000001?????????????????: sa = 5'd17;
            32'b0000000000000001????????????????: sa = 5'd16;
            32'b00000000000000001???????????????: sa = 5'd15;
            32'b000000000000000001??????????????: sa = 5'd14;
            32'b0000000000000000001?????????????: sa = 5'd13;
            32'b00000000000000000001????????????: sa = 5'd12;
            32'b000000000000000000001???????????: sa = 5'd11;
            32'b0000000000000000000001??????????: sa = 5'd10;
            32'b00000000000000000000001?????????: sa = 5'd9;
            32'b000000000000000000000001????????: sa = 5'd8;
            32'b0000000000000000000000001???????: sa = 5'd7;
            32'b00000000000000000000000001??????: sa = 5'd6;
            32'b000000000000000000000000001?????: sa = 5'd5;
            32'b0000000000000000000000000001????: sa = 5'd4;
            32'b00000000000000000000000000001???: sa = 5'd3;
            32'b000000000000000000000000000001??: sa = 5'd2;
            32'b0000000000000000000000000000001?: sa = 5'd1;
            default: sa = 5'd0;
        endcase
        tSig = i_unsigned[30:0] << (30 - sa);     //Normalized sig
        //Rounding to nearest (Ties To Even)
        if (tSig[6:0] > 7'b011_1111) begin        //Add 1 to the remaining bits
            roSig = tSig[30:7] + 1;
        end 
        else if (tSig[6:0] < 7'b011_1111) begin   //Do nothing
            roSig = tSig[30:7];
        end
        else begin                                //Check for tSig[7]: EVEN or ODD
            roSig = tSig[30:7] + tSig[7];
        end
        fExp =  i_unsigned ? (127 + sa + roSig[24]) : 8'b0;
    end
    assign f = {i[31] , fExp , roSig[22:0]};
endmodule